package shared_pkg;
	class shared;
		/*The signal will be defined as well as the 
		error_count and correct_count in a shared package that you will create named shared_pkg. */
		static int test_finished = 0;
		static int error_count   = 0;
		static int correct_count = 0;
	endclass
endpackage  